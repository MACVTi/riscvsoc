`include "./definitions.vh"

module cpu #(parameter VECTOR_RESET=32'h00000000, VECTOR_INTERRUPT = 32'h00000000) (


    );
endmodule
