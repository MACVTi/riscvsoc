// Written by Jack McEllin - 15170144
// Definitions for the immediate generator module

`ifndef _immgen_h_
    `define _immgen_h_

    //------------------------------------------------------------
	// ALU function select values
	//------------------------------------------------------------

	`define IMM_ITYPE	   3'b000		
    `define IMM_STYPE	   3'b001
    `define IMM_BTYPE	   3'b010
    `define IMM_UTYPE	   3'b011
    `define IMM_JTYPE	   3'b100
    `define IMM_RTYPE	   3'b101
    
`endif