// Written by Jack McEllin - 15170144
// Definitions for the load generator module

`ifndef _loadgen_h_
    `define _loadgen_h_

    //------------------------------------------------------------
	// Load generator select values
	//------------------------------------------------------------

	`define LOAD_LB    	   3'b000		
    `define LOAD_LH	       3'b001
    `define LOAD_LW	       3'b010
    `define LOAD_LBU	   3'b011
    `define LOAD_LHU	   3'b100
    
`endif