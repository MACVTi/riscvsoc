`ifndef _alu_h_
    `define _alu_h_

    //------------------------------------------------------------
	// Functions
	//------------------------------------------------------------

	`define ALU_ADD		   4'b0000		//ADD
	`define ALU_SUB		   4'b0001		//SUB
	`define ALU_SLL		   4'b0010		//SUB
	`define ALU_SLT		   4'b0011		//SUB
	`define ALU_SLTU       4'b0100		//SUB
	`define ALU_XOR		   4'b0101		//SUB
	`define ALU_SRL		   4'b0110		//SUB
	`define ALU_SRA	       4'b0111		//SUB
	`define ALU_OR		   4'b1000		//SUB
	`define ALU_AND        4'b1001		//SUB

`endif