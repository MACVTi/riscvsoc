// Written by Jack McEllin - 15170144
// Definitions for the store generator module

`ifndef _storegen_h_
    `define _storegen_h_

    //------------------------------------------------------------
	// Load generator select values
	//------------------------------------------------------------

	`define STORE_SB       3'b00		
    `define STORE_SH       3'b01
    `define STORE_SW       3'b10
    
`endif